module alu(
    input a,
    input b,
    input [2:0] op,
    output reg [7:0] out,
    output reg carry
);
    always_comb begin
        case (op)
            
        endcase
    end
endmodule
