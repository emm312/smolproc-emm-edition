module execute(
    input [7:0] op_a,
    input [7:0] op_b,
    input [7:0] opcode,
    input [7:0] dst,

    output reg [7:0] res
);

endmodule